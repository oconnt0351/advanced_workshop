/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_oconnt_counter (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // Internal register: 8-bit counter
  reg [7:0] count;

  // Sequential logic: counter increments on every clock
  always @(posedge clk) begin
    if (!rst_n)        // Active-low reset
      count <= 8'b0;
    else
      count <= count + 1;
  end

  // Assign counter to output
  assign uo_out = count;

  // Tie off unused IOs
  assign uio_out = 0;
  assign uio_oe  = 0;

  // Prevent warnings for unused signals
  wire _unused = &{ena, ui_in, uio_in, 1'b0};

endmodule
